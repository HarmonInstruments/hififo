`include "buildtime.vh"
`define USE_GT_DRP
`define NLANES 4
`define ENABLE 8'b01110111
